`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:05:34 05/14/2015 
// Design Name: 
// Module Name:    median5x5 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module median5x5 # (
	parameter [9:0] H_SIZE = 83
)(
		input binary,
		input de,
		input vsync,
		input hsync,
		
		output median
    );


endmodule
